//area of rectangle
module ex15;
integer l=10,w=5,f;
initial begin
f=(l*w);
$display("The area of rectangle is :%f",f);
end
endmodule

