//perform the given data's
module ex6(a,b,c,d,o0,o1,o2,o3,o4,o5,o6,o7);
input [3:0]a,b,c,d;
output [3:0]o0,o1,o2,o3,o4,o5,o6,o7 ;
assign o0=a|b;
assign o1=c&d;
assign o2=a^b;
assign o3=~(c^d);
assign o4=(c&&d);
assign o5=a||b;
assign o6=b>>2;
assign o7=a<<3;
endmodule

module tb;
reg [3:0]a,b,c,d;
wire [3:0]o0,o1,o2,o3,o4,o5,o6,o7;
ex6 i1(a,b,c,d,o0,o1,o2,o3,o4,o5,o6,o7);
initial begin
$monitor(" \n(a|b)=%b \n(c&d)=%b \n(a^b)=%b \n~(c^d)=%b \n(c&&d)=%b \n(a||b)=%b \n(b>>2)=%b \n(a<<3)=%b \n",o0,o1,o2,o3,o4,o5,o6,o7);
 a=7;b=4'b1001;c=4'hc;d=14;
end 
endmodule


