module x;
real x;
initial begin
x=198.12300000;
$display("Integer x=%d",x);
$display("Real x=%f",x);
end
endmodule
