module ex10;
reg [7:0]a=170,b=31,c=171,d=255;
initial begin
$monitor("%h,%h,%h,%h",a,b,c,d);
end 
endmodule
