//area of circle
module ex16;
integer r=2,f;
initial begin
f=2*(3.145*(r*r));
$display("The area of circle is :%f",f);
end
endmodule
