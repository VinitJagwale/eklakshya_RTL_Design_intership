module hi;
 initial 
  begin
  $display ("hello world verilog");
  $display ("hello world verilog");
  #10 $finish;
  end
endmodule

