module ex9;
reg [1:0]a=3,b=2,c=1,d=0;
initial begin 
$display("%b",a);
$display("%b",b);
$display("%b",c);
$display("%b",d);
$finish;
end
endmodule
