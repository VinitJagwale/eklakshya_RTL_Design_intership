module ex17;
real a=15,b=15.55,f;
initial begin
f=a*b;
$display("In Integer F= %d\nIn Real    F= %f",f,f);
end
endmodule 

